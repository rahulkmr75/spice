** modelling 741 op-amp **

*model transistrors
.MODEL Q741PNP PNP(IS=2E-15 RB=300 RC=300 RE=10 
+BF=50 BR=4 VA=50 TF=30NS CJE=.3PF PE=.55V ME=.5
+CJC=2PF PC=.55V MC=.5 CCS=3PF PS=.52V MS=.5V)

.MODEL SPNP PNP(IS=1E-14 RB=150 RC=50 RE=2 
+BR=4 BF=50 VA=50 TF=20NS CJE=.5PF PE=.55V ME=.5
+CJC=2PF PC=.52V MC=.5 CCS=3PF PS=.52V MS=.5V)

.MODEL Q741NPN NPN(IS=5E-15 RB=200 RC=250 BF=250 
+BR=2 RE=2 VA=130 TF=.35NS CJE=1PF PE=.7V ME=.33
+CJC=.3PF PC=.55V MC=.5 CCS=3PF PS=.52 MS=.5V)
*

*uA741 Operational Amp Spice File
.subckt lm_741_op_amp 1 2 20 Vcc=15V Vee=-15V
    *** 1= V+  , 2=V- 20=Vout ***
    ** 741 OP AMP **
    * BIAS CIRCUIT *
    Q12 23 23 21 Q741PNP
    Q11 24 24 22 Q741NPN
    Q10 6 24 26 Q741NPN
    Q13A 17 23 21 Q741PNP 1
    Q13B 14 23 21 Q741PNP 3
    Q15 17 18 20 Q741NPN
    Q21 25 19 20 Q741PNP
    Q22 8 25 22 Q741NPN
    Q24 25 25 22 Q741NPN
    Q23B 22 14 8 Q741PNP
    R5 23 24 39K
    R4 26 22 5K
    R11 25 22 50K
    CC 14 8 30PF
    *
    * DIFF AMP *
    Q1 3 1 4 Q741NPN
    Q2 3 2 5 Q741NPN
    Q3 7 6 4 Q741PNP
    Q4 8 6 5 Q741PNP
    Q5 7 9 10 Q741NPN
    Q6 8 9 11 Q741NPN
    Q7 21 7 9 Q741NPN
    Q8 3 3 21 Q741PNP
    Q9 6 3 21 Q741PNP
    R1 10 22 1K
    R2 11 22 1K
    R3 9 22 50K

    * DARLINGTON **
    Q16 21 8 12 Q741NPN
    Q17 14 12 13 Q741NPN
    R9 12 22 50K
    R8 13 22 100
    * OUTPUT STAGE *
    Q19 17 17 16 Q741NPN
    Q18 17 16 15 Q741NPN
    Q23A 22 14 15 Q741PNP
    Q14 21 17 18 Q741NPN 3
    Q20 22 15 19 SPNP
    R10 16 15 40K
    R6 18 20 27
    R7 20 19 22
    * POWER SUPPLY *
    VCC 21 0 DC= { Vcc}
    VEE 22 0 DC= {-Vcc}
.ends lm_741_op_amp
*

